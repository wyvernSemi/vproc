###################################################################
# Makefile for Virtual Processor VHDL testcode in Modelsim
#
# Copyright (c) 2005-2024 Simon Southwell.
#
# This file is part of VProc.
#
# VProc is free software: you can redistribute it and/or modify
# it under the terms of the GNU General Public License as published by
# the Free Software Foundation, either version 3 of the License, or
# (at your option) any later version.
#
# VProc is distributed in the hope that it will be useful,
# but WITHOUT ANY WARRANTY; without even the implied warranty of
# MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
# GNU General Public License for more details.
#
# You should have received a copy of the GNU General Public License
# along with VProc. If not, see <http://www.gnu.org/licenses/>.
#
###################################################################

###################################################################
# THIS FILE IS DEPRECATED AND IS FOR BACKWARDS COMPATIBILITY      #
###################################################################

# User overridable variables
HDL                = VHDL
USRFLAGS           =
OPTFLAG            = -g
USER_C             = VUserMain0.c VUserMain1.cpp
USRCDIR            = usercode
TESTDIR            = .
MEMC               =
MEMMODELDIR        = .

# Set up the common make command for the ModelSim/Questa makefile
COMMONCMD = $(MAKE) --no-print-directory            \
                    HDL="$(HDL)"                    \
                    USRFLAGS="$(USRFLAGS)"          \
                    OPTFLAG="$(OPTFLAG)"            \
                    USER_C="$(USER_C)"              \
                    USRCDIR="$(USRCDIR)"            \
                    TESTDIR="$(TESTDIR)"            \
                    MEMC="$(MEMC)"                  \
                    MEMMODELDIR="$(MEMMODELDIR)"    \
                    -f makefile

#------------------------------------------------------
# BUILD RULES
#------------------------------------------------------

all:
	@$(COMMONCMD)

#------------------------------------------------------
# EXECUTION RULES
#------------------------------------------------------

sim:
	@$(COMMONCMD) sim

run:
	@$(COMMONCMD) run

rungui:
	@$(COMMONCMD) rungui

gui: rungui

help:
	@$(COMMONCMD) help

clean:
	@$(COMMONCMD) clean
